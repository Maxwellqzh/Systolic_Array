`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Create Date:   2025/11/24
// Design Name:   PE_core
// Module Name:   PE_core
// Description:   ���ڼ�������8λ�з�������ˣ������봫�ݸ���һ����Ԫ�����ۼӽ��
// input:
//      clk: ʱ���ź�
//      rst_n: ��λ�ź�
//      a_curr: ��ǰ�����Aֵ
//      b_curr: ��ǰ�����Bֵ
// output:
//      a_last: ���ݸ���һ����Ԫ��Aֵ
//      b_last: ���ݸ���һ����Ԫ��Bֵ
//      data_out: �ۼӽ��
//

module PE_Core
#(parameter DATA_WIDTH = 8)
(
    input clk,rst_n,
    input signed [DATA_WIDTH-1:0] a_curr,
    input signed [DATA_WIDTH-1:0] b_curr,
    output reg signed [DATA_WIDTH-1:0] a_last,
    output reg signed [DATA_WIDTH-1:0] b_last,
    output reg signed [2*DATA_WIDTH-1:0] data_out
    );
    wire signed [2*DATA_WIDTH-1:0] data_tmp;
    wire rst;
    assign rst = !rst_n;
    always@(posedge clk or negedge rst_n)
        begin
            if(!rst_n)
                begin
                    a_last<='d0;
                    b_last<='d0;
                    data_out<='d0;
                end
            else
                begin
                    a_last<=a_curr;
                    b_last<=b_curr;
                    data_out<=data_out+data_tmp;
                end
        end

    // multiplier u_multiplier(
    //     .clk(clk),
    //     .CE(1),
    //     .SCLR(rst),
    //     .A(a_curr),
    //     .B(b_curr),
    //     .P (data_tmp)
    // );
    multiplier u_multiplier(
        .clk(clk),
        .CE(1),
        .SCLR(rst),
        .A(a_curr),
        .B(b_curr),
        .P(data_tmp)
    );
endmodule

module multiplier
#(parameter DATA_WIDTH = 8)
(
    input clk,CE,SCLR,
    input signed [DATA_WIDTH-1:0] A,
    input signed [DATA_WIDTH-1:0] B,
    output reg   [2*DATA_WIDTH-1:0] P
);
    always@(posedge clk or posedge SCLR)
        begin
            if(SCLR)
                P<=0;
            else
            if(CE)
                P<=A*B;
            else
                P<=P;
        end
endmodule
