// Engineer:      Zhenhang Qin
// Create Date:   2025/11/24
// Design Name:   PE_array
// Module Name:   PE_array
// Description:   ���ڼ�������������ˣ�������������֧��os��wsģʽ
// input:
//      clk: ʱ���ź�
//      rst_n: ��λ�ź�
//      en: �ⲿ����ʹ��
//      data_flow: ������ģʽѡ���ź�,1ΪWSģʽ,0ΪOSģʽ
//      load: Ȩ�ؼ���ʹ���ź�,��loadΪ1ʱ����B��ΪȨ������
//      acc_en: �ۼ�ʹ���ź�,��acc_enΪ1ʱ����C_acc��Ϊ�ۼ�����
//      A: �����Aֵ,����ΪROWS*DATA_WIDTH
//      B: �����Bֵ,����ΪCOLS*DATA_WIDTH
//      C_acc: �����C_accֵ,����ΪCOLS*2*DATA_WIDTH��������Ҫ����ˮ��ʽ����
// output:
//      valid: �����Ч�źţ���en����֮�󣬼��������֮�󣬵ȴ�������ɺ��Զ����߲����֣�ֱ�����н���������������
//      C_out: ������,�������,����ΪCOLS*2*DATA_WIDTH������WSģʽ��C_Out��Ҫ�ⲿ����

`timescale 1ns / 1ps

module PE_Array #(
    parameter DATA_WIDTH = 8,
    parameter ROWS = 8,
    parameter COLS = 8
)(
    input clk,
    input rst_n,
    input en,            // �ⲿ����ʹ��
    
    // --- �����ź� ---
    input data_flow,     // 1: WS Mode, 0: OS Mode
    input load,          // WS Weight Loading
    input acc_en,        // [����] �ۼ�ʹ��: 1=�ۼ�C_acc, 0=��0��ʼ���� (����WS����ģʽ��Ч)
    
    // --- �������� ---
    input signed [ROWS*DATA_WIDTH-1:0] A,
    input signed [COLS*DATA_WIDTH-1:0] B,
    input signed [COLS*2*DATA_WIDTH-1:0] C_acc,

    // --- ������� ---
    output valid,        // ���ڲ� Controller ����
    output signed [COLS*2*DATA_WIDTH-1:0] C_out, // ԭʼ��б����� (Raw Skewed Output)
);

    // =========================================================
    // 1. �ڲ����߶���
    // =========================================================
    wire signed [DATA_WIDTH-1:0] w_hor [0:ROWS-1][0:COLS];
    wire signed [2*DATA_WIDTH-1:0] w_ver [0:ROWS][0:COLS-1];
    
    // �ڲ������ź�
    wire internal_drain; 

    // =========================================================
    // 2. ʵ����״̬������
    // =========================================================
    PE_Status_Controller #(
        .ROWS(ROWS),
        .COLS(COLS)
    ) u_controller (
        .clk(clk),
        .rst_n(rst_n),
        .en(en),
        .data_flow(data_flow),
        .drain_out(internal_drain), // OSģʽʹ�õ� Drain �ź�
        .valid_out(valid)           // ȫ�������Ч�ź�
    );

    // =========================================================
    // 3. �߽����봦�� (�� Loopback Mux)
    // =========================================================
    genvar i, j;
    generate
        // --- ������� A ---
        for (i = 0; i < ROWS; i = i + 1) begin : A_Input_Map
            assign w_hor[i][0] = A[((i+1)*DATA_WIDTH)-1 -: DATA_WIDTH];
        end

        // --- �������� B / C_acc / 0 ---
        for (j = 0; j < COLS; j = j + 1) begin : B_Input_Map
            // ��ȡ��ǰ�е� B ���� (8-bit)
            wire signed [DATA_WIDTH-1:0] b_curr_col;
            assign b_curr_col = B[((j+1)*DATA_WIDTH)-1 -: DATA_WIDTH];
            
            // ��ȡ��ǰ�е� Loopback ���� (16-bit)
            wire signed [2*DATA_WIDTH-1:0] acc_curr_col;
            assign acc_curr_col = C_acc[((j+1)*2*DATA_WIDTH)-1 -: 2*DATA_WIDTH];

            // ��չ B �� 16-bit (������չ)
            wire signed [2*DATA_WIDTH-1:0] b_extended;
            assign b_extended = {{DATA_WIDTH{b_curr_col[DATA_WIDTH-1]}}, b_curr_col};

            // ����ѡ���߼���
            // 1. WS Load: ����ιȨ�� (B)
            // 2. OS Mode: ����ι������ (B)
            // 3. WS Compute & Acc_En: ι Loopback ���� (C_acc)
            // 4. WS Compute & !Acc_En: ι 0 (��ʼ��һ�ּ���)
            
            assign w_ver[0][j] = (data_flow && load) ? b_extended :   // WS: ����Ȩ��
                                 (!data_flow)        ? b_extended :   // OS: ������
                                 (acc_en)            ? acc_curr_col : // WS: �ۼӾɽ��
                                                       {(2*DATA_WIDTH){1'b0}}; // WS: �¼��� (����0)
        end
    endgenerate

    // =========================================================
    // 4. PE ��������
    // =========================================================
    generate
        for (i = 0; i < ROWS; i = i + 1) begin : Row_Gen
            for (j = 0; j < COLS; j = j + 1) begin : Col_Gen
                PE_Core #(
                    .DATA_WIDTH(DATA_WIDTH)
                ) u_pe (
                    .clk(clk),
                    .rst_n(rst_n),
                    .data_flow(data_flow),
                    .load(load),
                    .drain(internal_drain), 
                    
                    .left (w_hor[i][j]),       
                    .up   (w_ver[i][j]),       
                    .right(w_hor[i][j+1]),     
                    .down (w_ver[i+1][j])      
                );
            end
        end
    endgenerate

    // =========================================================
    // 5. �߽�������� 
    // =========================================================
    // ֱ��������еײ������ݣ�����б��ʱ���Ա��ⲿ Loopback ֱ�ӶԽ�
    generate
        for (j = 0; j < COLS; j = j + 1) begin : Final_Output_Map
            assign C_out[((j+1)*2*DATA_WIDTH)-1 -: 2*DATA_WIDTH] = w_ver[ROWS][j];
        end

        // A ͸�����
        for (i = 0; i < ROWS; i = i + 1) begin : A_Pass_Map
            assign A_pass_out[((i+1)*DATA_WIDTH)-1 -: DATA_WIDTH] = w_hor[i][COLS];
        end
    endgenerate

endmodule