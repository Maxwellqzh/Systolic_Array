// Engineer:      Zhenhang Qin
// Create Date:   2025/11/24
// Design Name:   PE_array
// Module Name:   PE_array
// Description:   ���ڼ�������������ˣ�����������
// input:
//      clk: ʱ���ź�
//      rst_n: ��λ�ź�
//      en: ����ʹ���ź�,�����һ�����ݵĵ�һ��Ԫ�������ʹ������
//      A: �����Aֵ,����ΪROWS*DATA_WIDTH
//      B: �����Bֵ,����ΪCOLS*DATA_WIDTH
//      C: ������,�������
//      valid: �����Ч�źţ�������ɺ�����һ��ʱ������

`timescale 1ns / 1ps


module PE_Array #(
    parameter DATA_WIDTH = 8,
    parameter ROWS = 8,
    parameter COLS = 8
)(
    input clk,
    input rst_n,
    
    // --- �����ź� (���ⲿ Controller �ṩ) ---
    input data_flow,     // 1: WS Mode, 0: OS Mode
    input load,          // WS Weight Loading
    input drain,         // OS Result Draining
    
    // --- �������� ---
    // A (Left Input): ÿһ��һ�� 8-bit ����
    input signed [ROWS*DATA_WIDTH-1:0] A,

    // B (Top Input): ÿһ��һ�� 8-bit ����
    input signed [COLS*DATA_WIDTH-1:0] B,

    // --- ������� ---
    // C (Bottom Output): ÿһ��һ�� 16-bit ���
    // ע�⣺����Ǵӵײ�����ˮ��һ���������ģ��������������������
    output signed [COLS*2*DATA_WIDTH-1:0] C_out,
    
    // ����/�����ã����Ҳ�� A ��� (��ѡ)
    output signed [ROWS*DATA_WIDTH-1:0] A_pass_out
);

    // =========================================================
    // 1. �ڲ����߶��� (Interconnects)
    // =========================================================
    // ˮƽ���� (Horizontal Wires): ���� A
    // �ߴ�: [ROWS] �� x [COLS+1] �� (��������������������)
    wire signed [DATA_WIDTH-1:0] w_hor [0:ROWS-1][0:COLS];

    // ��ֱ���� (Vertical Wires): ���� B / Partial Sum / Result
    // �ߴ�: [ROWS+1] �� x [COLS] �� (����������������)
    // ע��λ���� 2*DATA_WIDTH (16-bit)
    wire signed [2*DATA_WIDTH-1:0] w_ver [0:ROWS][0:COLS-1];

    // =========================================================
    // 2. �߽����봦�� (Boundary Inputs)
    // =========================================================
    
    genvar i, j;
    generate
        // --- ������� A ---
        for (i = 0; i < ROWS; i = i + 1) begin : A_Input_Map
            assign w_hor[i][0] = A[((i+1)*DATA_WIDTH)-1 -: DATA_WIDTH];
        end

        // --- �������� B / Partial Sum ---
        for (j = 0; j < COLS; j = j + 1) begin : B_Input_Map
            wire signed [DATA_WIDTH-1:0] b_curr_col;
            assign b_curr_col = B[((j+1)*DATA_WIDTH)-1 -: DATA_WIDTH];

            // �߼�ѡ��
            // Case 1: WS����ģʽ (data_flow=1, load=0) -> ��������� 0 (���ֺͳ�ʼֵ)
            // Case 2: ������� (WS���� / OSģʽ) -> ������ B (��չ��16λ)
            // ע�������չ (Sign Extension)
            
            assign w_ver[0][j] = (data_flow && !load) ? 
                                 {(2*DATA_WIDTH){1'b0}} :  // WS����: ι0
                                 {{DATA_WIDTH{b_curr_col[DATA_WIDTH-1]}}, b_curr_col}; // ����: ιB (������չ)
        end
    endgenerate

    // =========================================================
    // 3. PE �������� (Array Instantiation)
    // =========================================================
    generate
        for (i = 0; i < ROWS; i = i + 1) begin : Row_Gen
            for (j = 0; j < COLS; j = j + 1) begin : Col_Gen
                
                PE_Core #(
                    .DATA_WIDTH(DATA_WIDTH)
                ) u_pe (
                    .clk(clk),
                    .rst_n(rst_n),
                    
                    // �����źŹ㲥
                    .data_flow(data_flow),
                    .load(load),
                    .drain(drain),
                    
                    // ��������
                    .left (w_hor[i][j]),       // �������
                    .up   (w_ver[i][j]),       // ��������
                    .right(w_hor[i][j+1]),     // �����ұ�
                    .down (w_ver[i+1][j])      // ��������
                );
                
            end
        end
    endgenerate

    // =========================================================
    // 4. �߽�������� (Boundary Outputs)
    // =========================================================
    generate
        // --- �ײ���� (Result / Drain) ---
        // ȡ�� w_ver �����һ��
        for (j = 0; j < COLS; j = j + 1) begin : C_Output_Map
            assign C_out[((j+1)*2*DATA_WIDTH)-1 -: 2*DATA_WIDTH] = w_ver[ROWS][j];
        end

        // --- �Ҳ���� (A͸����ͨ�����ڵ��Ի���) ---
        for (i = 0; i < ROWS; i = i + 1) begin : A_Pass_Map
            assign A_pass_out[((i+1)*DATA_WIDTH)-1 -: DATA_WIDTH] = w_hor[i][COLS];
        end
    endgenerate

endmodule