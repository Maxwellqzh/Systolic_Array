// Engineer:      Zhenhang Qin
// Create Date:   2025/11/24
// Design Name:   PE_core
// Module Name:   PE_Core
// Description:   ���ڼ�������8λ�з�������ˣ������봫�ݸ���һ����Ԫ�����ۼӽ����֧��WS��OS����ģʽ
// input:
//      clk: ʱ���ź�
//      rst_n: ��λ�ź�'
//      drain: ������ʹ���ź�,�ߵ�ƽʱOS״̬��������
//      data_flow: ģʽѡ���źţ�1ΪWSģʽ��0ΪOSģʽ
//      load: Ȩ�ؼ���ʹ���ź�,�ߵ�ƽʱ��data_in������ΪȨ������
//      left: ˮƽ����A
//      up: ��ֱ���룬Loadģʽ��ΪȨ�أ�����ģʽ��Ϊ�Ϸ�������Partial Sum
// output:
//      right: ˮƽ���A
//      down: ��ֱ�����Loadģʽ�´���Ȩ�أ�����ģʽ������ۼӽ��

`timescale 1ns / 1ps

module PE_Core #(
    parameter DATA_WIDTH = 8
)(
    input clk,
    input rst_n,
    input data_flow,            // 1: WS, 0: OS
    input load,                 // WSģʽ����Ȩ��
    input drain,                // OSģʽ������ʹ��
    input signed [DATA_WIDTH-1:0] left,      
    input signed [2*DATA_WIDTH-1:0] up,  
    
    output reg signed [DATA_WIDTH-1:0] right,     
    output reg signed [2*DATA_WIDTH-1:0] down
);

    reg signed [DATA_WIDTH-1:0] weight_reg; 
    reg signed [2*DATA_WIDTH-1:0] ps_reg;   
    reg drain_1d;
    wire drain_neg;
    wire signed [2*DATA_WIDTH-1:0] temp_result;

    // ����ʵ�ʽ���˷���B�˿ڵ��ź�
    // WSģʽ: �ñ��ش�õ� weight_reg
    // OSģʽ: ֱ������������ up (��ȡ��8λ)������1���ӳ�
    wire signed [DATA_WIDTH-1:0] mult_input_b;
    assign mult_input_b = (data_flow) ? weight_reg : up[DATA_WIDTH-1:0];

    // ʵ�����˷���
    multiplier u_multiplier(
        .clk(clk),
        .CE(1'b1),
        .SCLR(!rst_n),
        .A(left),
        .B(mult_input_b), // ʹ��ѡ�����ź�
        .P(temp_result)
    );

    always@(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            drain_1d <= 0;
        end else begin
            drain_1d <= drain;
        end
    end

    assign drain_neg = drain_1d && !drain;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            right      <= 0;
            down       <= 0;
            weight_reg <= 0;
            ps_reg     <= 0;
        end else begin
            // 1. ˮƽ����͸�� (��������ģʽ)
            right <= left;

            if (data_flow) begin
                // ========================
                // WS Mode (Weight Stationary)
                // ========================
                if (load) begin
                    // Ȩ�ؼ����봫��
                    weight_reg <= up[DATA_WIDTH-1:0];
                    down       <= up;
                end else begin
                    // Ȩ�ز��������ֺ�����
                    // down = �Ϸ��Ĳ��ֺ� + ��ǰ�˻�
                    down <= up + temp_result;
                end
            end else begin
                // ========================
                // OS Mode (Output Stationary)
                // ========================
                // Ȩ�ر������� (���ݸ��·�PE)
                down <= up; 
                if (drain || drain_1d) begin
                    // ����ģʽ��ֹͣ�ۼӣ������ͨ�� down �³�ȥ
                    // ��ʱ down �������������������ٴ�Ȩ��
                    // ���drain�����һ�����ڣ������������ɣ����м��ۼ�����
                    if(drain_1d)
                        down <= up; 
                    else
                        down <= ps_reg; 
                    if(drain_neg)      
                        ps_reg <= 0;
                    else
                        ps_reg <= ps_reg;
                end else begin
                    // �ۼ�ģʽ
                    ps_reg <= ps_reg + temp_result;
                end
            end
        end
    end
endmodule

module multiplier
#(parameter DATA_WIDTH = 8)
(
    input clk,CE,SCLR,
    input signed [DATA_WIDTH-1:0] A,
    input signed [DATA_WIDTH-1:0] B,
    output reg   [2*DATA_WIDTH-1:0] P
);
    always@(posedge clk or posedge SCLR)
        begin
            if(SCLR)
                P<=0;
            else
            if(CE)
                P<=A*B;
            else
                P<=P;
        end
endmodule
