// Engineer:      Zhenhang Qin
// Create Date:   2025/11/24
// Design Name:   PE_array
// Module Name:   PE_array
// Description:   ���ڼ�������������ˣ�����������
// input:
//      clk: ʱ���ź�
//      rst_n: ��λ�ź�
//      en: ����ʹ���ź�,�����һ�����ݵĵ�һ��Ԫ�������ʹ������
//      A: �����Aֵ,����ΪROWS*DATA_WIDTH
//      B: �����Bֵ,����ΪCOLS*DATA_WIDTH
//      C: ������,�������
//      valid: �����Ч�źţ�������ɺ�����һ��ʱ������

`timescale 1ns / 1ps


module PE_Array #(
    parameter DATA_WIDTH = 8,
    parameter ROWS = 8,
    parameter COLS = 8
)(
    input clk,
    input rst_n,
    input en,  // ����ʹ���ź�,�����һ�����������ʹ������

    // ������� A���������룩��չƽΪһά����
    // ���з�ʽ��A[0], A[1], ..., A[ROWS-1]
    input signed [ROWS*DATA_WIDTH-1:0] A,

    // �������� B���������룩��չƽΪһά����  
    // ���з�ʽ��B[0], B[1], ..., B[COLS-1]
    input signed [COLS*DATA_WIDTH-1:0] B,

    // ������� C���ۼӣ���չƽΪһά����
    // ���з�ʽ��C[0][0], C[0][1], ..., C[0][COLS-1], C[1][0], ...
    output signed [ROWS*COLS*2*DATA_WIDTH-1:0] C,
    
    output valid  // �����Ч�ź�
);

// �ڲ������ź�
wire signed [DATA_WIDTH-1:0] A_2d [0:ROWS-1];
wire signed [DATA_WIDTH-1:0] B_2d [0:COLS-1];
wire signed [2*DATA_WIDTH-1:0] C_2d [0:ROWS-1][0:COLS-1];

// PE֮��������ź�
wire signed [DATA_WIDTH-1:0] a_horizontal [0:ROWS-1][0:COLS];  // ˮƽ���򴫲���A����
wire signed [DATA_WIDTH-1:0] b_vertical   [0:ROWS][0:COLS-1];  // ��ֱ���򴫲���B����

// ��ˮ�߿����ź�
reg [ROWS+COLS-1:0] pipeline_valid;  // ��ˮ����Ч��־
wire computation_done;  // ��������ź�

// ������ˮ����ȣ����ݴ����뵽�����Ҫ��ʱ�䣩
localparam PIPELINE_DEPTH = ROWS + COLS - 1;

// ������Aչƽ����ά����
genvar i, j;
generate
    for (i = 0; i < ROWS; i = i + 1) begin : A_reshape
        assign A_2d[i] = A[(i+1)*DATA_WIDTH-1 : i*DATA_WIDTH];
    end
    
    // ������Bչƽ����ά����  
    for (i = 0; i < COLS; i = i + 1) begin : B_reshape
        assign B_2d[i] = B[(i+1)*DATA_WIDTH-1 : i*DATA_WIDTH];
    end
    
    // �������뵽PE���б߽�
    for (i = 0; i < ROWS; i = i + 1) begin : A_input_conn
        assign a_horizontal[i][0] = A_2d[i];  // ÿ�еĵ�һ��PE�����ⲿA����
    end
    
    for (j = 0; j < COLS; j = j + 1) begin : B_input_conn
        assign b_vertical[0][j] = B_2d[j];    // ÿ�еĵ�һ��PE�����ⲿB����
    end
    
    // ����PE����
    for (i = 0; i < ROWS; i = i + 1) begin : row_gen
        for (j = 0; j < COLS; j = j + 1) begin : col_gen
            PE_Core #(
                .DATA_WIDTH(DATA_WIDTH)
            ) PE_inst (
                .clk(clk),
                .rst_n(rst_n),
                .a_curr(a_horizontal[i][j]),      // ��ǰPE��A����
                .b_curr(b_vertical[i][j]),        // ��ǰPE��B����
                .a_last(a_horizontal[i][j+1]),    // A������Ҳ�PE
                .b_last(b_vertical[i+1][j]),      // B������·�PE
                .data_out(C_2d[i][j])             // ���������
            );
            
        end
    end
    
    // �����C_2dչƽ��һά�������
    for (i = 0; i < ROWS; i = i + 1) begin : C_output_row
        for (j = 0; j < COLS; j = j + 1) begin : C_output_col
            assign C[((i*COLS + j) + 1) * (2*DATA_WIDTH) - 1 : 
                     (i*COLS + j) * (2*DATA_WIDTH)] = C_2d[i][j];
        end
    end
    
endgenerate

// �����Ч�źţ����������������ʹ���Ѿ����ͣ���ʾ�������һ�����ݣ�
reg en_delayed;
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        en_delayed <= 0;
    end else begin
        en_delayed <= en;
    end
end

// ���en���½��أ��Ӹߵ��ͣ�
wire en_falling_edge = en_delayed && !en;

// ��ˮ����Ч��־����
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        pipeline_valid <= 0;
    end else begin
        // ��λ�Ĵ�����������������ˮ���е�λ��
        pipeline_valid <= {pipeline_valid[ROWS+COLS-2:0], en_falling_edge};
    end
end

// ��������жϣ������һ��PE��������Чʱ�������������
assign computation_done = pipeline_valid[PIPELINE_DEPTH-1];


// ��Ч�ź����ɣ�����⵽en�½��غ󣬵ȴ��������
reg valid_generation;
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        valid_generation <= 0;
    end else if (en_falling_edge) begin
        // ��⵽en�½��أ���ʼ�ȴ��������
        valid_generation <= 1;
    end else if (computation_done && valid_generation) begin
        // ������ɣ������Ч���ɱ�־
        valid_generation <= 0;
    end
end

// ������Ч�ź����
assign valid = computation_done && valid_generation;

endmodule