`timescale 1ns / 1ps

module tb_Systolic_input_controller;

    // ��������
    parameter DATA_WIDTH = 8;
    parameter ROWS = 4;
    parameter COLS = 4;
    parameter CLK_PERIOD = 10;

    // �źŶ���
    reg clk;
    reg rst_n;
    reg enable;
    reg signed [DATA_WIDTH*ROWS-1:0] A;
    reg signed [DATA_WIDTH*COLS-1:0] B;
    wire signed [DATA_WIDTH*ROWS-1:0] A_out;
    wire signed [DATA_WIDTH*COLS-1:0] B_out;
    wire valid;

    // ��������������������鿴��
    reg [DATA_WIDTH-1:0] A_in_array [0:ROWS-1];
    reg [DATA_WIDTH-1:0] B_in_array [0:COLS-1];
    reg [DATA_WIDTH-1:0] A_out_array [0:ROWS-1];
    reg [DATA_WIDTH-1:0] B_out_array [0:COLS-1];

    // ��ʱ�������
    reg [DATA_WIDTH-1:0] temp_A [0:ROWS-1];
    reg [DATA_WIDTH-1:0] temp_B [0:COLS-1];

    // ʵ��������ģ��
    Systolic_input_controller #(
        .DATA_WIDTH(DATA_WIDTH),
        .ROWS(ROWS),
        .COLS(COLS)
    ) uut (
        .clk(clk),
        .rst_n(rst_n),
        .enable(enable),
        .A(A),
        .B(B),
        .A_out(A_out),
        .B_out(B_out),
        .valid(valid)
    );

    // ʱ������
    always #(CLK_PERIOD/2) clk = ~clk;

    // ���񣺽��������ת��Ϊ����
    task update_output_arrays;
        integer i;
        begin
            for (i = 0; i < ROWS; i = i + 1) begin
                A_out_array[i] = A_out[((i+1)*DATA_WIDTH)-1 -: DATA_WIDTH];
            end
            for (i = 0; i < COLS; i = i + 1) begin
                B_out_array[i] = B_out[((i+1)*DATA_WIDTH)-1 -: DATA_WIDTH];
            end
        end
    endtask

    // ����������������
    task set_input_data_A;
        input [DATA_WIDTH-1:0] a0, a1, a2, a3;
        integer i;
        begin
            temp_A[0] = a0;
            temp_A[1] = a1;
            temp_A[2] = a2;
            temp_A[3] = a3;
            
            for (i = 0; i < ROWS; i = i + 1) begin
                A_in_array[i] = temp_A[i];
                A[((i+1)*DATA_WIDTH)-1 -: DATA_WIDTH] = temp_A[i];
            end
        end
    endtask

    task set_input_data_B;
        input [DATA_WIDTH-1:0] b0, b1, b2, b3;
        integer i;
        begin
            temp_B[0] = b0;
            temp_B[1] = b1;
            temp_B[2] = b2;
            temp_B[3] = b3;
            
            for (i = 0; i < COLS; i = i + 1) begin
                B_in_array[i] = temp_B[i];
                B[((i+1)*DATA_WIDTH)-1 -: DATA_WIDTH] = temp_B[i];
            end
        end
    endtask

    // ������ʾ�����������
    task display_arrays;
        integer i;
        begin
            $write("����: A_in_array = [");
            for (i = 0; i < ROWS; i = i + 1) begin
                $write("%0d", A_in_array[i]);
                if (i < ROWS-1) $write(", ");
            end
            $write("]");
            
            $write("  B_in_array = [");
            for (i = 0; i < COLS; i = i + 1) begin
                $write("%0d", B_in_array[i]);
                if (i < COLS-1) $write(", ");
            end
            $write("]\n");
            
            $write("���: A_out_array = [");
            for (i = 0; i < ROWS; i = i + 1) begin
                $write("%0d", A_out_array[i]);
                if (i < ROWS-1) $write(", ");
            end
            $write("]");
            
            $write("  B_out_array = [");
            for (i = 0; i < COLS; i = i + 1) begin
                $write("%0d", B_out_array[i]);
                if (i < COLS-1) $write(", ");
            end
            $write("]");
            
            $display("  valid = %0d", valid);
        end
    endtask

    // ������
    initial begin
        // ��ʼ��
        clk = 0;
        rst_n = 0;
        enable = 0;
        A = 0;
        B = 0;

        // ��ʼ������
        for (integer i = 0; i < ROWS; i = i + 1) begin
            A_in_array[i] = 0;
            A_out_array[i] = 0;
            temp_A[i] = 0;
        end
        for (integer i = 0; i < COLS; i = i + 1) begin
            B_in_array[i] = 0;
            B_out_array[i] = 0;
            temp_B[i] = 0;
        end

        // ��λ
        #(CLK_PERIOD * 2);
        rst_n = 1;
        #(CLK_PERIOD);

        $display("=== Starting Test ===");
        $display("Testing enable high for 4 cycles, input different A, B data each cycle");

        // �׶�1: enable����4�����ڣ�ÿ���������벻ͬ����
        $display("\n--- Phase 1: enable high for 4 cycles, input different data ---");
        enable = 1;
        
        // ����1: �����һ������
        set_input_data_A(1, 2, 3, 4);
        set_input_data_B(5, 6, 7, 8);
        #(CLK_PERIOD);
        update_output_arrays();
        $display("Cycle 1:");
        display_arrays();
        
        // ����2: ����ڶ�������
        set_input_data_A(10, 20, 30, 40);
        set_input_data_B(50, 60, 70, 80);
        #(CLK_PERIOD);
        update_output_arrays();
        $display("Cycle 2:");
        display_arrays();
        
        // ����3: �������������
        set_input_data_A(100, 200, 300, 400);
        set_input_data_B(500, 600, 700, 800);
        #(CLK_PERIOD);
        update_output_arrays();
        $display("Cycle 3:");
        display_arrays();
        
        // ����4: �������������
        set_input_data_A(11, 22, 33, 44);
        set_input_data_B(55, 66, 77, 88);
        #(CLK_PERIOD);
        update_output_arrays();
        $display("Cycle 4:");
        display_arrays();

        // �׶�2: enable����3�����ڣ��۲���λЧ��
        $display("\n--- Phase 2: enable low for 3 cycles, observe shifting ---");
        enable = 0;
        
        // ��������
        set_input_data_A(0, 0, 0, 0);
        set_input_data_B(0, 0, 0, 0);
        
        #(CLK_PERIOD);
        update_output_arrays();
        $display("Cycle 5:");
        display_arrays();
        
        #(CLK_PERIOD);
        update_output_arrays();
        $display("Cycle 6:");
        display_arrays();
        
        #(CLK_PERIOD);
        update_output_arrays();
        $display("Cycle 7:");
        display_arrays();

        $display("\n=== Test Finished ===");
        #(CLK_PERIOD * 2);
        $finish;
    end

    // ���μ�¼
    initial begin
        $dumpfile("tb_Systolic_input_controller.vcd");
        $dumpvars(0, tb_Systolic_input_controller);
    end

endmodule