// Engineer:      Zhenhang Qin
// Create Date:   2025/11/24
// Design Name:   controller
// Module Name:   controller
// Description:   �������������źţ������������A��B�źŷ�ʱ����
// input:
//      clk: ʱ���ź�
//      rst_n: ��λ�ź�
//      enable: ����ʹ���ź�,�����һ���������������
//      A: �����Aֵ,����ΪROWS*DATA_WIDTH
//      B: �����Bֵ,����ΪCOLS*DATA_WIDTH
// output:
//      valid: enable���ӳ��źţ����ڿ���PE_array������ʹ���ź�

module Systolic_Input_Controller #(
    parameter DATA_WIDTH = 8,
    parameter ROWS = 8,
    parameter COLS = 8
)(
    input clk,
    input rst_n, 
    input enable,
    input signed [DATA_WIDTH*ROWS-1:0] A,  // չƽ��A����
    input signed [DATA_WIDTH*COLS-1:0] B,  // չƽ��B����
    output signed [DATA_WIDTH*ROWS-1:0] A_out,
    output signed [DATA_WIDTH*COLS-1:0] B_out,
    output reg valid
);

    // A����λ�Ĵ����飨ÿ��һ����
    reg signed [DATA_WIDTH-1:0] A_shift [0:ROWS-1][0:ROWS-1];
    // B����λ�Ĵ����飨ÿ��һ����  
    reg signed [DATA_WIDTH-1:0] B_shift [0:COLS-1][0:COLS-1];
    
    integer i, j, k, m;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            valid <= 0;
        end
        else if (enable) begin
            valid <= 1;
        end
        else begin
            valid <= 0;
        end
    end
    
    // ��ʼ����λ�Ĵ���
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            for (i = 0; i < ROWS; i = i + 1) begin
                for (j = 0; j < ROWS; j = j + 1) begin
                    A_shift[i][j] <= 0;
                end
            end
            for (i = 0; i < COLS; i = i + 1) begin
                for (j = 0; j < COLS; j = j + 1) begin
                    B_shift[i][j] <= 0;
                end
            end
        end
        else begin
            // A������λ�߼�
            for (i = 0; i < ROWS; i = i + 1) begin
                for (j = 0; j < i; j = j + 1) begin
                    A_shift[i][j] <= A_shift[i][j+1];
                end
                // ��Verilog�Ĳ���ѡ���﷨
                A_shift[i][i] <= A[((i+1)*DATA_WIDTH)-1 -: DATA_WIDTH];
            end
            
            // B������λ�߼�
            for (i = 0; i < COLS; i = i + 1) begin
                for (j = 0; j < i; j = j + 1) begin
                    B_shift[i][j] <= B_shift[i][j+1];
                end
                // ��Verilog�Ĳ���ѡ���﷨
                B_shift[i][i] <= B[((i+1)*DATA_WIDTH)-1 -: DATA_WIDTH];
            end
        end
    end
    
    // �����ǰ�Խ�������
    genvar gi, gj;
    generate
        for (gi = 0; gi < ROWS; gi = gi + 1) begin : A_OUTPUT_GEN
            assign A_out[((gi+1)*DATA_WIDTH)-1 -: DATA_WIDTH] = A_shift[gi][0];
        end
        for (gj = 0; gj < COLS; gj = gj + 1) begin : B_OUTPUT_GEN
            assign B_out[((gj+1)*DATA_WIDTH)-1 -: DATA_WIDTH] = B_shift[gj][0];
        end
    endgenerate

endmodule